`timescale 1ns / 1ps
`include "nroot.v"


module nroot_tb;
   wire [31:0]result;
    wire underflow,overflow;

    reg [31:0]	A;
	reg	[31:0]	B;
	reg			CLK,RST;


    nroot uut(	.A(A),
                .B(B),
				.CLK(CLK),
				.RST(RST),
                .overflow(overflow),
                .underflow(underflow),
                .result(result));

always
begin
#0	CLK = 1'B0;
#2	CLK = 1'B1;
#2;
end

initial
        begin
	/////////////////////////////////////////////////////////////////////
	
			A = 32'b01001100111100000101001101110000; //1.26E8
			B = 32'b01000010111101100000000000000000; //123
			#1 RST = 1'B1;
			#5 RST = 1'B0;
			#5 RST = 1'B1;
			#12000;
			
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b00111100101111100000110111101101; //0.232
//	        	B = 32'b01000001010010101011100001010010; //12.67
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//			
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b01000010000100001100001010001111; //36.19
//			B = 32'b00111111001000111101011100001010; //0.64
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b00111111010001100110011001100110; //0.775
//	        	B = 32'b00111111001010111000010100011111; //0.67
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//
//	/////////////////////////////////////////////////////////////////////
//
//			A = 32'b00111110100000000000000000000000; //0.25
//			B = 32'b10111110100000110110111000101111; //-0.2567
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b00000000000000000000000000000000; //0
//			B = 32'b00000000000000000000000000000000; //0
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b01111111100000000000000000000000; //Inf
//			B = 32'b00000000000000000000000000000000; //0
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//			
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b00000000000000000000000000000000; //0
//			B = 32'b01111111100000000000000000000000; //Inf
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//			
//	///////////////////////////////////////////////////////////////////	
//
//			A = 32'b01111111100000000000000000000000; //Inf
//			B = 32'b01111111100000000000000000000000; //Inf
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//			
//	/////////////////////////////////////////////////////////////////////
//	
//			A = 32'b01111111100000000000000000000000; //Inf
//			B = 32'b11111111111111111111111111111111; //NaN
//			#1 RST = 1'B1;
//			#5 RST = 1'B0;
//			#5 RST = 1'B1;
//			#12000;
//			
//	/////////////////////////////////////////////////////////////////////		
			$finish;
        end
		
initial
begin
$vcdplusfile("tb_nroot.vpd");
$vcdpluson();
end

endmodule
