
module MUL_wallace_tree_24_tb( );
	
reg [24-1:0]in1,in2;
wire[49-1:0]out;

mul_wallace_tree_24 MUL_0(.in1(in1),.in2(in2),.out(out));
initial begin
	in1 = 24'h123456;

	in2 = 24'h852;
	#10;
	in1 = 24'h1;

	in2 = 24'h153;
	#10;
	in1 = 24'h945698;

	in2 = 24'h123549;
	#10;
	
	in1 = 24'h523321;

    in2 = 24'h851662;
    #10;
    in1 = 24'h7861;

    in2 = 24'h870153;
    #10;
    in1 = 24'h855781;

    in2 = 24'h123069;
    #10;
	in1 = 24'h523561;

    in2 = 24'h852352;
    #10;
    in1 = 24'h1235;

    in2 = 24'h168553;
    #10;
    in1 = 24'h809512;

    in2 = 24'h341239;
    #10;
    
	in1 = 24'h521255;

    in2 = 24'h852532;
    #10;
    in1 = 24'h12;

    in2 = 24'h15345;
    #10;
    in1 = 24'h812351;

    in2 = 24'h1239;
    #10;
	// in1 = 32'b01000000000000000000000000000000;

	// in2 = 32'b00111111100000000000000000000000;
	// #10;

	// in1 = 32'b01000000000000000000000000000000;

	// in2 = 32'b01000000000000000000000000000000;
	// #10;
	
	// in1 = 32'b01000000101010000000000000000000;

	// in2 = 32'b01000000000000000000000000000000;
	// #10;
	// in1 = 32'b10111111100000000000000000000000; //-1

	// in2 = 32'b01000000000000000000000000000000;
	// #10;
	// in1 = 32'b01000000001000000000000000000000; //2.5

	// in2 = 32'b01000000011000000000000000000000; //3.5
	// #10;
	// in1 = 32'b01000100111111000111001100110011; //2019.6
	
	// in2 = 32'b11000000011000000000000000000000; //-3.5
	// #10;

	// in1 = 32'b01000100111111000111001100110011; //2019.6
	
	// in2 = 32'b11111111100000000000000000000001;// NaN

	// #10;
	// in1 = 32'b0_00000000_00000000000000000000000; // 0
	
	// in2 = 32'b0_00000000_00000000000000000000000; // 0

	// #10;
	// in1 = 32'b1_11111111_00000000000000000000000;// -INF
	
	// in2 = 32'b0_11111111_00000000000000000000000;// +INF

	// #10;
	// in1 = 32'b0_11111111_00000000000000000000000;// +INF
	
	// in2 = 32'b0_00000000_00000000000000000000000;// 0

	// #10;
	// in1 = 32'b1_11111111_00000000000000000000000;// -INF
	
	// in2 = 32'b1_11111111_00000000000000000000000;// -INF

	// #10;
	// in1 = 32'b0_11111111_00000000000000000000000;// +INF
	
	// in2 = 32'b1_11111111_00000000000000000000000;// -INF



end
	
endmodule 