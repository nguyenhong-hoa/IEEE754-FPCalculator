module MUX_23_1(
	select,
	in,
	out
);

input [4:0] select;
input [31:0] in;
output out;




endmodule
